//=========================================================================
// Name & Email must be EXACTLY as in Gradescope roster!
// Name: Michelle Dozal
// Email: mdoza001@ucr.edu
//
// Assignment name: Lab #3 Pre-lab
// Lab section: 021
// TA: Yujia Zhai
//
// I hereby certify that I have not received assistance on this assignment,
// or used code, from ANY outside source other than the instruction team
// (apart from what was provided in the starter file).
//
//=========================================================================
`timescale 1ns/1ps

module datapath_tb;
    reg clk;
    reg[5:0] instr_op;
    reg[5:0] instr_field;
    reg[8:0] R;
    wire[8:0] result;
    wire[3:0] alu_result;
    reg[3:0] R_alu_result;
    
    //unit under test
    controlUnit uut(
        .instr_op(instr_op),
        .reg_dst(result[8]),
        .alu_src(result[7]),
        .mem_to_reg(result[6]),
        .reg_write(result[5]),
        .mem_read(result[4]),
        .mem_write(result[3]),
        .branch(result[2]),
        .alu_op(result[1:0])
    );
    
    aluControlUnit uut2(
        .alu_op(result[1:0]),
        .instruction_5_0(instr_field),
        .alu_out(alu_result)
);
    
    
    initial begin
    clk = 1;
    forever begin
    clk = ~clk; #50;
    end
    end

    integer failedTests = 0;
    integer totalTests = 0;

    initial begin
    //@(posedge clk);
    #10
    
        $write("Test Group 1: Testing Main Contol Unit... \n");
        $write("\tTest Case 1.1: R-format...");
        totalTests = totalTests + 1;
        instr_op = 6'b000000;
        R = 9'b100100010;
        #100;
        if(R !== result)begin
            $write("failed: expected: %b, got %b\n", R, result);
            failedTests = failedTests + 1;
        end else begin
            $write("passed\n");
        end

        $write("\tTest Case 1.2: lw...");
        totalTests = totalTests + 1;
        instr_op = 6'b100011;
        R = 9'b011110000;
        #100;
        if(R !== result) begin
           $write("failed: expected: %b, got %b\n", R, result);
           failedTests = failedTests + 1;
        end else begin
           $write("passed\n");
        end
        #10;

        
        totalTests = totalTests + 1;
        $write("\tTest Case 1.3: sw...");
        instr_op = 6'b101011;
        R = 9'bx1x001000;
        #100;
        if (R !== result) begin
            $write("failed: expected: %b, got %b\n", R, result);
            failedTests  = failedTests + 1;
        end else begin
            $write("passed\n");
        end
        #10;
        
        totalTests = totalTests + 1;
        $write("\tTest Case 1.4: beq...");
        instr_op = 6'b000100;
        R = 9'bx0x000101;
        #100;
        if (R !== result) begin
            $write("failed: expected: %b, got %b\n", R, result);
            failedTests  = failedTests + 1;
        end else begin
            $write("passed\n");
        end
        #10;

        totalTests = totalTests + 1;
        $write("\tTest Case 1.5: addi,subi...");
        instr_op = 6'b001000;
        R = 9'b110100010;
        #100;
        if (R !== result) begin
            $write("failed: expected: %b, got %b\n", R, result);
            failedTests  = failedTests + 1;
        end else begin
            $write("passed\n");
        end
        #10;
        
        totalTests = totalTests + 1;
        $write("Test Group 2: ALU...\n");
        $write("\tTest Case 2.1: R-type opcode add...");
        instr_op = 6'b000000;
        // alu_op will be generated by controlUnit.v
        instr_field = 6'b100000;
        R_alu_result = 4'b0010;
        #100;
        if (R_alu_result !== alu_result) begin
            $write("failed: expected: %b, got %b\n", R_alu_result, alu_result);
            failedTests  = failedTests + 1;
        end else begin
            $write("passed\n");
        end
        #10;

        totalTests = totalTests + 1;
        $write("\tTest Case 2.2: R-type opcode sub...");
        instr_op = 6'b000000;
        // alu_op will be generated by controlUnit.v
        instr_field = 6'b100010;
        R_alu_result = 4'b0110;
        #100;
        if (R_alu_result !== alu_result) begin
            $write("failed: expected: %b, got %b\n", R_alu_result, alu_result);
            failedTests  = failedTests + 1;
        end else begin
            $write("passed\n");
        end
        #10
        
        totalTests = totalTests + 1;
        $write("\tTest Case 2.3: R-type opcode AND...");
        instr_op = 6'b000000;
        // alu_op will be generated by controlUnit.v
        instr_field = 6'b100100;
        R_alu_result = 4'b0000;
        #100;
        if (R_alu_result !== alu_result) begin
            $write("failed: expected: %b, got %b\n", R_alu_result, alu_result);
            failedTests  = failedTests + 1;
        end else begin
            $write("passed\n");
        end
        #10;

        totalTests = totalTests + 1;
        $write("\tTest Case 2.4: R-type opcode OR...");
        instr_op = 6'b000000;
        // alu_op will be generated by controlUnit.v
        instr_field = 6'b100101;
        R_alu_result = 4'b0001;
        #100;
        if (R_alu_result !== alu_result) begin
            $write("failed: expected: %b, got %b\n", R_alu_result, alu_result);
            failedTests  = failedTests + 1;
        end else begin
            $write("passed\n");
        end
        #10;

        totalTests = totalTests + 1;
        $write("\tTest Case 2.5: R-type opcode NOR...");
        instr_op = 6'b000000;
        // alu_op will be generated by controlUnit.v
        instr_field = 6'b100111;
        R_alu_result = 4'b1100;
        #100;
        if (R_alu_result !== alu_result) begin
            $write("failed: expected: %b, got %b\n", R_alu_result, alu_result);
            failedTests  = failedTests + 1;
        end else begin
            $write("passed\n");
        end
        #10;

        totalTests = totalTests + 1;
        $write("\tTest Case 2.6: R-type opcode SLT...");
        instr_op = 6'b000000;
        // alu_op will be generated by controlUnit.v
        instr_field = 6'b101010;
        R_alu_result = 4'b0111;
        #100;
        if (R_alu_result !== alu_result) begin
            $write("failed: expected: %b, got %b\n", R_alu_result, alu_result);
            failedTests  = failedTests + 1;
        end else begin
            $write("passed\n");
        end
        #10;

        $write("\n--------------------------------------------------------------");
        $write("\nTesting complete\nPassed %0d / %0d tests",totalTests-failedTests,totalTests);
        $write("\n--------------------------------------------------------------\n");
        $finish();

end

endmodule
